`include "decoder.svh"

module decoder(
    input logic [31:0] inst_i,
    input logic fetch_err_i,
    output is_t is_o
);

    always_comb begin
        unique casez(inst_i)
            32'b010011??????????????????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_LI;
                is_o.alu_op = `_ALU_STYPE_PCPLUS4;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd1;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = `_FUSEL_EX_ALU;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S16;
                is_o.branch_type = `_BRANCH_NOCONDITION;
                is_o.target_type = `_TARGET_ABS;
                is_o.cmp_type = 3'd0;
            end
            32'b010100??????????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd1;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = `_FUSEL_EX_ALU;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = `_BRANCH_NOCONDITION;
                is_o.target_type = `_TARGET_REL;
                is_o.cmp_type = 3'd0;
            end
            32'b010101??????????????????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_LI;
                is_o.alu_op = `_ALU_STYPE_PCPLUS4;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd1;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = `_FUSEL_EX_ALU;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_BL1;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = `_BRANCH_NOCONDITION;
                is_o.target_type = `_TARGET_REL;
                is_o.cmp_type = 3'd0;
            end
            32'b010110??????????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd1;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd1;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RD;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S16;
                is_o.branch_type = `_BRANCH_CONDITION;
                is_o.target_type = `_TARGET_REL;
                is_o.cmp_type = `_CMP_E;
            end
            32'b010111??????????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd1;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd1;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RD;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S16;
                is_o.branch_type = `_BRANCH_CONDITION;
                is_o.target_type = `_TARGET_REL;
                is_o.cmp_type = `_CMP_NE;
            end
            32'b011000??????????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd1;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd1;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RD;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S16;
                is_o.branch_type = `_BRANCH_CONDITION;
                is_o.target_type = `_TARGET_REL;
                is_o.cmp_type = `_CMP_LT;
            end
            32'b011001??????????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd1;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd1;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RD;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S16;
                is_o.branch_type = `_BRANCH_CONDITION;
                is_o.target_type = `_TARGET_REL;
                is_o.cmp_type = `_CMP_GE;
            end
            32'b011010??????????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd1;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd1;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RD;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S16;
                is_o.branch_type = `_BRANCH_CONDITION;
                is_o.target_type = `_TARGET_REL;
                is_o.cmp_type = `_CMP_LTU;
            end
            32'b011011??????????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd1;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd1;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RD;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S16;
                is_o.branch_type = `_BRANCH_CONDITION;
                is_o.target_type = `_TARGET_REL;
                is_o.cmp_type = `_CMP_GEU;
            end
            32'b0001010?????????????????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_LI;
                is_o.alu_op = `_ALU_STYPE_LUI;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd1;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = `_FUSEL_EX_ALU;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_IMM;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_S20;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0001110?????????????????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_LI;
                is_o.alu_op = `_ALU_STYPE_PCADDUI;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd1;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = `_FUSEL_EX_ALU;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_IMM;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_S20;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000100????????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd1;
                is_o.refetch = 1'd1;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd1;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd1;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd1;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd1;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = `_FUSEL_M2_CSR;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RD;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00100000????????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = `_MEM_TYPE_WORD;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd1;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd1;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd1;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S14;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00100001????????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = `_MEM_TYPE_WORD;
                is_o.mem_write = 1'd1;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd1;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd1;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RD;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S14;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0000001000??????????????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_CMP;
                is_o.alu_op = `_ALU_STYPE_SLT;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd1;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd1;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_IMM;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_S12;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0000001001??????????????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_CMP;
                is_o.alu_op = `_ALU_STYPE_SLTU;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd1;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd1;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_IMM;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_S12;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0000001010??????????????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_INT;
                is_o.alu_op = `_ALU_STYPE_ADD;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd1;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd1;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_IMM;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_S12;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0000001101??????????????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_BW;
                is_o.alu_op = `_ALU_STYPE_AND;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd1;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = `_FUSEL_EX_ALU;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_IMM;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U12;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0000001110??????????????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_BW;
                is_o.alu_op = `_ALU_STYPE_OR;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd1;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = `_FUSEL_EX_ALU;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_IMM;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U12;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0000001111??????????????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_BW;
                is_o.alu_op = `_ALU_STYPE_XOR;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd1;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = `_FUSEL_EX_ALU;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_IMM;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U12;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0000011000??????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd1;
                is_o.refetch = 1'd1;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = `_MEM_TYPE_BYTE;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd1;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd1;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S12;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0010100000??????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = `_MEM_TYPE_BYTE;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd1;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd1;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S12;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0010100001??????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = `_MEM_TYPE_HALF;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd1;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd1;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S12;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0010100010??????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = `_MEM_TYPE_WORD;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd1;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd1;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S12;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0010100100??????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = `_MEM_TYPE_BYTE;
                is_o.mem_write = 1'd1;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd1;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RD;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S12;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0010100101??????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = `_MEM_TYPE_HALF;
                is_o.mem_write = 1'd1;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd1;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RD;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S12;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0010100110??????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = `_MEM_TYPE_WORD;
                is_o.mem_write = 1'd1;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd1;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RD;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S12;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0010101000??????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = `_MEM_TYPE_UBYTE;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd1;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd1;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S12;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0010101001??????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = `_MEM_TYPE_UHALF;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd1;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd1;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S12;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0010101011??????????????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000000100000???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_INT;
                is_o.alu_op = `_ALU_STYPE_ADD;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd1;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd1;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000000100010???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_INT;
                is_o.alu_op = `_ALU_STYPE_SUB;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd1;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd1;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000000100100???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_CMP;
                is_o.alu_op = `_ALU_STYPE_SLT;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd1;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd1;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000000100101???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_CMP;
                is_o.alu_op = `_ALU_STYPE_SLTU;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd1;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd1;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000000101000???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_BW;
                is_o.alu_op = `_ALU_STYPE_NOR;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd1;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = `_FUSEL_EX_ALU;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000000101001???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_BW;
                is_o.alu_op = `_ALU_STYPE_AND;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd1;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = `_FUSEL_EX_ALU;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000000101010???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_BW;
                is_o.alu_op = `_ALU_STYPE_OR;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd1;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = `_FUSEL_EX_ALU;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000000101011???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_BW;
                is_o.alu_op = `_ALU_STYPE_XOR;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd1;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = `_FUSEL_EX_ALU;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000000101110???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_SFT;
                is_o.alu_op = `_ALU_STYPE_SLL;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd1;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000000101111???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_SFT;
                is_o.alu_op = `_ALU_STYPE_SRL;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd1;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000000110000???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_SFT;
                is_o.alu_op = `_ALU_STYPE_SRA;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd1;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000000111000???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_MUL;
                is_o.alu_op = `_MUL_TYPE_MULL;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd1;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd1;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000000111001???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_MUL;
                is_o.alu_op = `_MUL_TYPE_MULH;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd1;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd1;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000000111010???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_MUL;
                is_o.alu_op = `_MUL_TYPE_MULHU;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd1;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd1;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000001000000???????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = `_DIV_TYPE_DIV;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd1;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd1;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = `_FUSEL_WB_DIV;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000001000001???????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = `_DIV_TYPE_MOD;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd1;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd1;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = `_FUSEL_WB_DIV;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000001000010???????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = `_DIV_TYPE_DIVU;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd1;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd1;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = `_FUSEL_WB_DIV;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000001000011???????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = `_DIV_TYPE_MODU;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd1;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd1;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd1;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = `_FUSEL_WB_DIV;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000001010110???????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd1;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000001010110???????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd1;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd1;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000010000001???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_SFT;
                is_o.alu_op = `_ALU_STYPE_SLL;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd1;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_IMM;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000010001001???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_SFT;
                is_o.alu_op = `_ALU_STYPE_SRL;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd1;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_IMM;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000000010010001???????????????: begin
                is_o.alu_grand_op = `_ALU_GTYPE_SFT;
                is_o.alu_op = `_ALU_STYPE_SRA;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd1;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = `_FUSEL_M1_ALU;
                is_o.fu_sel_m2 = `_FUSEL_M2_ALU;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_IMM;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_RD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000110010010001???????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd1;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd1;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd1;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00000110010010011???????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd1;
                is_o.refetch = 1'd1;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd1;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd1;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd1;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd1;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_RK;
                is_o.reg_type_r1 = `_REG_R1_RJ;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00111000011100100???????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd1;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b00111000011100101???????????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd1;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd1;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0000000000000000011000??????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = `_RDCNT_ID_VLOW;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd1;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd1;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = `_FUSEL_M2_CSR;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R0_NONE;
                is_o.reg_type_w = `_REG_W_RJD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0000000000000000011001??????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = `_RDCNT_VHIGH;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd1;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = `_FUSEL_M2_CSR;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_RJD;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0000011001001000001010??????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd1;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd1;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd1;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0000011001001000001011??????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd1;
                is_o.refetch = 1'd1;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd1;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd1;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0000011001001000001100??????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd1;
                is_o.refetch = 1'd1;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd1;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd1;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0000011001001000001101??????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd1;
                is_o.refetch = 1'd1;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd1;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd1;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            32'b0000011001001000001110??????????: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd1;
                is_o.priv_inst = 1'd1;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = inst_i;
                is_o.need_csr = 1'd1;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = `_REG_R0_NONE;
                is_o.reg_type_r1 = `_REG_R1_NONE;
                is_o.reg_type_w = `_REG_W_NONE;
                is_o.imm_type = `_IMM_U5;
                is_o.addr_imm_type = `_ADDR_IMM_S26;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
            default: begin
                is_o.alu_grand_op = 2'd0;
                is_o.alu_op = 2'd0;
                is_o.ertn_inst = 1'd0;
                is_o.priv_inst = 1'd0;
                is_o.refetch = 1'd0;
                is_o.wait_inst = 1'd0;
                is_o.invalid_inst = 1'd0;
                is_o.syscall_inst = 1'd0;
                is_o.break_inst = 1'd0;
                is_o.csr_op_en = 1'd0;
                is_o.csr_rdcnt = 2'd0;
                is_o.tlbsrch_en = 1'd0;
                is_o.tlbrd_en = 1'd0;
                is_o.tlbwr_en = 1'd0;
                is_o.tlbfill_en = 1'd0;
                is_o.invtlb_en = 1'd0;
                is_o.mem_type = 3'd0;
                is_o.mem_write = 1'd0;
                is_o.mem_read = 1'd0;
                is_o.mem_cacop = 1'd0;
                is_o.llsc_inst = 1'd0;
                is_o.ibarrier = 1'd0;
                is_o.dbarrier = 1'd0;
                is_o.debug_inst = 32'd0;
                is_o.need_csr = 1'd0;
                is_o.need_mul = 1'd0;
                is_o.need_div = 1'd0;
                is_o.need_lsu = 1'd0;
                is_o.need_bpu = 1'd0;
                is_o.latest_r0_ex = 1'd0;
                is_o.latest_r0_m1 = 1'd0;
                is_o.latest_r0_m2 = 1'd0;
                is_o.latest_r0_wb = 1'd0;
                is_o.latest_r1_ex = 1'd0;
                is_o.latest_r1_m1 = 1'd0;
                is_o.latest_r1_m2 = 1'd0;
                is_o.latest_r1_wb = 1'd0;
                is_o.fu_sel_ex = 1'd0;
                is_o.fu_sel_m1 = 2'd0;
                is_o.fu_sel_m2 = 2'd0;
                is_o.fu_sel_wb = 1'd0;
                is_o.reg_type_r0 = 2'd0;
                is_o.reg_type_r1 = 1'd0;
                is_o.reg_type_w = 2'd0;
                is_o.imm_type = 3'd0;
                is_o.addr_imm_type = 2'd0;
                is_o.branch_type = 2'd0;
                is_o.target_type = 1'd0;
                is_o.cmp_type = 3'd0;
            end
        endcase
    end

endmodule
