`timescale 1ns/1ps
`ifndef _COMMON_HEADER
`define _COMMON_HEADER

// `define _DIFFTEST_ENABLE
`define _VERILATOR
// `define _FPGA
// `define _LUT_REG
// `define _ASIC

`define _CACHE_BUS_DATA_LEN (32)
`define _AXI_BURST_SIZE (4'b0011)
`define _SIMPLIFY_MUL (1)    // 0 for using multiplier 

`endif
