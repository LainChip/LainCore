// Generator : SpinalHDL v1.9.2    git head : 457a28dd4b2ae1f3a1f3ef4268c3a7f613ec81ed
// Component : decoder
// Git hash  : 2410ee731f2c9a14f8bfeec9a0ac79cf1bbe9426

`timescale 1ns/1ps

module decoder (
  input      [31:0]   inst_i,
  input               fetch_err_i,
  output     [95:0]   is_o
);

  wire       [31:0]   _zz_ctrl;
  wire       [31:0]   _zz_ctrl_1;
  wire                _zz_ctrl_2;
  wire       [0:0]    _zz_ctrl_3;
  wire                _zz_ctrl_4;
  wire       [31:0]   _zz_ctrl_5;
  wire       [0:0]    _zz_ctrl_6;
  wire       [31:0]   _zz_ctrl_7;
  wire       [31:0]   _zz_ctrl_8;
  wire       [53:0]   _zz_ctrl_9;
  wire                _zz_ctrl_10;
  wire       [0:0]    _zz_ctrl_11;
  wire                _zz_ctrl_12;
  wire       [31:0]   _zz_ctrl_13;
  wire       [0:0]    _zz_ctrl_14;
  wire       [31:0]   _zz_ctrl_15;
  wire       [31:0]   _zz_ctrl_16;
  wire       [49:0]   _zz_ctrl_17;
  wire                _zz_ctrl_18;
  wire       [0:0]    _zz_ctrl_19;
  wire                _zz_ctrl_20;
  wire       [31:0]   _zz_ctrl_21;
  wire       [31:0]   _zz_ctrl_22;
  wire                _zz_ctrl_23;
  wire       [31:0]   _zz_ctrl_24;
  wire       [0:0]    _zz_ctrl_25;
  wire       [31:0]   _zz_ctrl_26;
  wire       [31:0]   _zz_ctrl_27;
  wire       [1:0]    _zz_ctrl_28;
  wire                _zz_ctrl_29;
  wire       [31:0]   _zz_ctrl_30;
  wire                _zz_ctrl_31;
  wire       [31:0]   _zz_ctrl_32;
  wire       [0:0]    _zz_ctrl_33;
  wire                _zz_ctrl_34;
  wire       [31:0]   _zz_ctrl_35;
  wire       [0:0]    _zz_ctrl_36;
  wire       [31:0]   _zz_ctrl_37;
  wire       [31:0]   _zz_ctrl_38;
  wire       [1:0]    _zz_ctrl_39;
  wire                _zz_ctrl_40;
  wire       [31:0]   _zz_ctrl_41;
  wire                _zz_ctrl_42;
  wire       [31:0]   _zz_ctrl_43;
  wire       [45:0]   _zz_ctrl_44;
  wire                _zz_ctrl_45;
  wire       [31:0]   _zz_ctrl_46;
  wire       [0:0]    _zz_ctrl_47;
  wire       [31:0]   _zz_ctrl_48;
  wire       [31:0]   _zz_ctrl_49;
  wire                _zz_ctrl_50;
  wire                _zz_ctrl_51;
  wire       [31:0]   _zz_ctrl_52;
  wire       [0:0]    _zz_ctrl_53;
  wire       [2:0]    _zz_ctrl_54;
  wire                _zz_ctrl_55;
  wire       [0:0]    _zz_ctrl_56;
  wire       [31:0]   _zz_ctrl_57;
  wire       [0:0]    _zz_ctrl_58;
  wire       [31:0]   _zz_ctrl_59;
  wire       [41:0]   _zz_ctrl_60;
  wire                _zz_ctrl_61;
  wire       [0:0]    _zz_ctrl_62;
  wire       [31:0]   _zz_ctrl_63;
  wire       [1:0]    _zz_ctrl_64;
  wire       [31:0]   _zz_ctrl_65;
  wire       [31:0]   _zz_ctrl_66;
  wire       [31:0]   _zz_ctrl_67;
  wire       [31:0]   _zz_ctrl_68;
  wire       [0:0]    _zz_ctrl_69;
  wire       [1:0]    _zz_ctrl_70;
  wire       [31:0]   _zz_ctrl_71;
  wire       [31:0]   _zz_ctrl_72;
  wire       [31:0]   _zz_ctrl_73;
  wire       [31:0]   _zz_ctrl_74;
  wire       [39:0]   _zz_ctrl_75;
  wire                _zz_ctrl_76;
  wire       [31:0]   _zz_ctrl_77;
  wire       [31:0]   _zz_ctrl_78;
  wire       [0:0]    _zz_ctrl_79;
  wire                _zz_ctrl_80;
  wire       [37:0]   _zz_ctrl_81;
  wire       [0:0]    _zz_ctrl_82;
  wire                _zz_ctrl_83;
  wire       [31:0]   _zz_ctrl_84;
  wire       [0:0]    _zz_ctrl_85;
  wire       [31:0]   _zz_ctrl_86;
  wire       [31:0]   _zz_ctrl_87;
  wire       [34:0]   _zz_ctrl_88;
  wire                _zz_ctrl_89;
  wire       [4:0]    _zz_ctrl_90;
  wire       [31:0]   _zz_ctrl_91;
  wire       [31:0]   _zz_ctrl_92;
  wire                _zz_ctrl_93;
  wire       [31:0]   _zz_ctrl_94;
  wire       [0:0]    _zz_ctrl_95;
  wire       [31:0]   _zz_ctrl_96;
  wire       [31:0]   _zz_ctrl_97;
  wire       [1:0]    _zz_ctrl_98;
  wire                _zz_ctrl_99;
  wire       [31:0]   _zz_ctrl_100;
  wire                _zz_ctrl_101;
  wire       [31:0]   _zz_ctrl_102;
  wire                _zz_ctrl_103;
  wire                _zz_ctrl_104;
  wire       [31:0]   _zz_ctrl_105;
  wire       [0:0]    _zz_ctrl_106;
  wire       [31:0]   _zz_ctrl_107;
  wire       [31:0]   _zz_ctrl_108;
  wire       [2:0]    _zz_ctrl_109;
  wire                _zz_ctrl_110;
  wire       [31:0]   _zz_ctrl_111;
  wire       [0:0]    _zz_ctrl_112;
  wire       [31:0]   _zz_ctrl_113;
  wire       [31:0]   _zz_ctrl_114;
  wire       [0:0]    _zz_ctrl_115;
  wire       [31:0]   _zz_ctrl_116;
  wire       [31:0]   _zz_ctrl_117;
  wire       [0:0]    _zz_ctrl_118;
  wire       [0:0]    _zz_ctrl_119;
  wire       [31:0]   _zz_ctrl_120;
  wire       [31:0]   _zz_ctrl_121;
  wire       [5:0]    _zz_ctrl_122;
  wire                _zz_ctrl_123;
  wire       [31:0]   _zz_ctrl_124;
  wire       [0:0]    _zz_ctrl_125;
  wire       [31:0]   _zz_ctrl_126;
  wire       [31:0]   _zz_ctrl_127;
  wire       [3:0]    _zz_ctrl_128;
  wire                _zz_ctrl_129;
  wire       [31:0]   _zz_ctrl_130;
  wire       [0:0]    _zz_ctrl_131;
  wire       [31:0]   _zz_ctrl_132;
  wire       [31:0]   _zz_ctrl_133;
  wire       [1:0]    _zz_ctrl_134;
  wire                _zz_ctrl_135;
  wire       [31:0]   _zz_ctrl_136;
  wire                _zz_ctrl_137;
  wire       [31:0]   _zz_ctrl_138;
  wire       [30:0]   _zz_ctrl_139;
  wire       [4:0]    _zz_ctrl_140;
  wire                _zz_ctrl_141;
  wire       [31:0]   _zz_ctrl_142;
  wire       [0:0]    _zz_ctrl_143;
  wire       [31:0]   _zz_ctrl_144;
  wire       [31:0]   _zz_ctrl_145;
  wire       [2:0]    _zz_ctrl_146;
  wire                _zz_ctrl_147;
  wire       [31:0]   _zz_ctrl_148;
  wire       [0:0]    _zz_ctrl_149;
  wire       [31:0]   _zz_ctrl_150;
  wire       [31:0]   _zz_ctrl_151;
  wire       [0:0]    _zz_ctrl_152;
  wire       [31:0]   _zz_ctrl_153;
  wire       [31:0]   _zz_ctrl_154;
  wire                _zz_ctrl_155;
  wire       [0:0]    _zz_ctrl_156;
  wire       [0:0]    _zz_ctrl_157;
  wire       [31:0]   _zz_ctrl_158;
  wire       [31:0]   _zz_ctrl_159;
  wire       [27:0]   _zz_ctrl_160;
  wire                _zz_ctrl_161;
  wire                _zz_ctrl_162;
  wire       [31:0]   _zz_ctrl_163;
  wire       [0:0]    _zz_ctrl_164;
  wire       [3:0]    _zz_ctrl_165;
  wire                _zz_ctrl_166;
  wire       [31:0]   _zz_ctrl_167;
  wire       [0:0]    _zz_ctrl_168;
  wire       [31:0]   _zz_ctrl_169;
  wire       [31:0]   _zz_ctrl_170;
  wire       [1:0]    _zz_ctrl_171;
  wire                _zz_ctrl_172;
  wire       [31:0]   _zz_ctrl_173;
  wire                _zz_ctrl_174;
  wire       [31:0]   _zz_ctrl_175;
  wire       [25:0]   _zz_ctrl_176;
  wire                _zz_ctrl_177;
  wire       [0:0]    _zz_ctrl_178;
  wire       [31:0]   _zz_ctrl_179;
  wire       [31:0]   _zz_ctrl_180;
  wire       [4:0]    _zz_ctrl_181;
  wire                _zz_ctrl_182;
  wire       [31:0]   _zz_ctrl_183;
  wire       [0:0]    _zz_ctrl_184;
  wire       [31:0]   _zz_ctrl_185;
  wire       [31:0]   _zz_ctrl_186;
  wire       [2:0]    _zz_ctrl_187;
  wire                _zz_ctrl_188;
  wire       [31:0]   _zz_ctrl_189;
  wire       [0:0]    _zz_ctrl_190;
  wire       [31:0]   _zz_ctrl_191;
  wire       [31:0]   _zz_ctrl_192;
  wire       [0:0]    _zz_ctrl_193;
  wire       [31:0]   _zz_ctrl_194;
  wire       [31:0]   _zz_ctrl_195;
  wire       [0:0]    _zz_ctrl_196;
  wire       [5:0]    _zz_ctrl_197;
  wire                _zz_ctrl_198;
  wire       [31:0]   _zz_ctrl_199;
  wire       [0:0]    _zz_ctrl_200;
  wire       [31:0]   _zz_ctrl_201;
  wire       [31:0]   _zz_ctrl_202;
  wire       [3:0]    _zz_ctrl_203;
  wire                _zz_ctrl_204;
  wire       [31:0]   _zz_ctrl_205;
  wire       [0:0]    _zz_ctrl_206;
  wire       [31:0]   _zz_ctrl_207;
  wire       [31:0]   _zz_ctrl_208;
  wire       [1:0]    _zz_ctrl_209;
  wire                _zz_ctrl_210;
  wire       [31:0]   _zz_ctrl_211;
  wire                _zz_ctrl_212;
  wire       [31:0]   _zz_ctrl_213;
  wire       [23:0]   _zz_ctrl_214;
  wire                _zz_ctrl_215;
  wire       [0:0]    _zz_ctrl_216;
  wire       [31:0]   _zz_ctrl_217;
  wire       [31:0]   _zz_ctrl_218;
  wire       [0:0]    _zz_ctrl_219;
  wire       [31:0]   _zz_ctrl_220;
  wire       [31:0]   _zz_ctrl_221;
  wire       [0:0]    _zz_ctrl_222;
  wire       [0:0]    _zz_ctrl_223;
  wire       [31:0]   _zz_ctrl_224;
  wire       [31:0]   _zz_ctrl_225;
  wire       [21:0]   _zz_ctrl_226;
  wire                _zz_ctrl_227;
  wire                _zz_ctrl_228;
  wire       [31:0]   _zz_ctrl_229;
  wire       [0:0]    _zz_ctrl_230;
  wire       [1:0]    _zz_ctrl_231;
  wire                _zz_ctrl_232;
  wire       [31:0]   _zz_ctrl_233;
  wire                _zz_ctrl_234;
  wire       [31:0]   _zz_ctrl_235;
  wire       [19:0]   _zz_ctrl_236;
  wire                _zz_ctrl_237;
  wire       [0:0]    _zz_ctrl_238;
  wire       [31:0]   _zz_ctrl_239;
  wire       [31:0]   _zz_ctrl_240;
  wire       [4:0]    _zz_ctrl_241;
  wire                _zz_ctrl_242;
  wire       [31:0]   _zz_ctrl_243;
  wire       [0:0]    _zz_ctrl_244;
  wire       [31:0]   _zz_ctrl_245;
  wire       [31:0]   _zz_ctrl_246;
  wire       [2:0]    _zz_ctrl_247;
  wire                _zz_ctrl_248;
  wire       [31:0]   _zz_ctrl_249;
  wire       [0:0]    _zz_ctrl_250;
  wire       [31:0]   _zz_ctrl_251;
  wire       [31:0]   _zz_ctrl_252;
  wire       [0:0]    _zz_ctrl_253;
  wire       [31:0]   _zz_ctrl_254;
  wire       [31:0]   _zz_ctrl_255;
  wire       [0:0]    _zz_ctrl_256;
  wire       [5:0]    _zz_ctrl_257;
  wire                _zz_ctrl_258;
  wire       [31:0]   _zz_ctrl_259;
  wire       [0:0]    _zz_ctrl_260;
  wire       [31:0]   _zz_ctrl_261;
  wire       [31:0]   _zz_ctrl_262;
  wire       [3:0]    _zz_ctrl_263;
  wire                _zz_ctrl_264;
  wire       [31:0]   _zz_ctrl_265;
  wire       [0:0]    _zz_ctrl_266;
  wire       [31:0]   _zz_ctrl_267;
  wire       [31:0]   _zz_ctrl_268;
  wire       [1:0]    _zz_ctrl_269;
  wire                _zz_ctrl_270;
  wire       [31:0]   _zz_ctrl_271;
  wire                _zz_ctrl_272;
  wire       [31:0]   _zz_ctrl_273;
  wire       [17:0]   _zz_ctrl_274;
  wire                _zz_ctrl_275;
  wire       [0:0]    _zz_ctrl_276;
  wire       [31:0]   _zz_ctrl_277;
  wire       [31:0]   _zz_ctrl_278;
  wire       [3:0]    _zz_ctrl_279;
  wire                _zz_ctrl_280;
  wire       [31:0]   _zz_ctrl_281;
  wire       [0:0]    _zz_ctrl_282;
  wire       [31:0]   _zz_ctrl_283;
  wire       [31:0]   _zz_ctrl_284;
  wire       [1:0]    _zz_ctrl_285;
  wire                _zz_ctrl_286;
  wire       [31:0]   _zz_ctrl_287;
  wire                _zz_ctrl_288;
  wire       [31:0]   _zz_ctrl_289;
  wire       [0:0]    _zz_ctrl_290;
  wire       [1:0]    _zz_ctrl_291;
  wire                _zz_ctrl_292;
  wire       [31:0]   _zz_ctrl_293;
  wire                _zz_ctrl_294;
  wire       [31:0]   _zz_ctrl_295;
  wire       [15:0]   _zz_ctrl_296;
  wire                _zz_ctrl_297;
  wire       [0:0]    _zz_ctrl_298;
  wire       [31:0]   _zz_ctrl_299;
  wire       [31:0]   _zz_ctrl_300;
  wire       [3:0]    _zz_ctrl_301;
  wire                _zz_ctrl_302;
  wire       [31:0]   _zz_ctrl_303;
  wire       [0:0]    _zz_ctrl_304;
  wire       [31:0]   _zz_ctrl_305;
  wire       [31:0]   _zz_ctrl_306;
  wire       [1:0]    _zz_ctrl_307;
  wire                _zz_ctrl_308;
  wire       [31:0]   _zz_ctrl_309;
  wire                _zz_ctrl_310;
  wire       [31:0]   _zz_ctrl_311;
  wire       [0:0]    _zz_ctrl_312;
  wire       [9:0]    _zz_ctrl_313;
  wire                _zz_ctrl_314;
  wire       [31:0]   _zz_ctrl_315;
  wire       [0:0]    _zz_ctrl_316;
  wire       [31:0]   _zz_ctrl_317;
  wire       [31:0]   _zz_ctrl_318;
  wire       [7:0]    _zz_ctrl_319;
  wire                _zz_ctrl_320;
  wire       [31:0]   _zz_ctrl_321;
  wire       [0:0]    _zz_ctrl_322;
  wire       [31:0]   _zz_ctrl_323;
  wire       [31:0]   _zz_ctrl_324;
  wire       [5:0]    _zz_ctrl_325;
  wire                _zz_ctrl_326;
  wire       [31:0]   _zz_ctrl_327;
  wire       [0:0]    _zz_ctrl_328;
  wire       [31:0]   _zz_ctrl_329;
  wire       [31:0]   _zz_ctrl_330;
  wire       [31:0]   _zz_ctrl_331;
  wire       [3:0]    _zz_ctrl_332;
  wire                _zz_ctrl_333;
  wire       [31:0]   _zz_ctrl_334;
  wire       [31:0]   _zz_ctrl_335;
  wire       [31:0]   _zz_ctrl_336;
  wire       [0:0]    _zz_ctrl_337;
  wire                _zz_ctrl_338;
  wire       [31:0]   _zz_ctrl_339;
  wire       [31:0]   _zz_ctrl_340;
  wire       [31:0]   _zz_ctrl_341;
  wire       [1:0]    _zz_ctrl_342;
  wire       [0:0]    _zz_ctrl_343;
  wire                _zz_ctrl_344;
  wire       [31:0]   _zz_ctrl_345;
  wire       [31:0]   _zz_ctrl_346;
  wire       [31:0]   _zz_ctrl_347;
  wire       [0:0]    _zz_ctrl_348;
  wire                _zz_ctrl_349;
  wire       [31:0]   _zz_ctrl_350;
  wire       [31:0]   _zz_ctrl_351;
  wire       [31:0]   _zz_ctrl_352;
  wire       [13:0]   _zz_ctrl_353;
  wire                _zz_ctrl_354;
  wire                _zz_ctrl_355;
  wire       [31:0]   _zz_ctrl_356;
  wire       [0:0]    _zz_ctrl_357;
  wire       [3:0]    _zz_ctrl_358;
  wire                _zz_ctrl_359;
  wire       [31:0]   _zz_ctrl_360;
  wire       [0:0]    _zz_ctrl_361;
  wire       [31:0]   _zz_ctrl_362;
  wire       [31:0]   _zz_ctrl_363;
  wire       [1:0]    _zz_ctrl_364;
  wire                _zz_ctrl_365;
  wire       [31:0]   _zz_ctrl_366;
  wire                _zz_ctrl_367;
  wire       [31:0]   _zz_ctrl_368;
  wire       [11:0]   _zz_ctrl_369;
  wire                _zz_ctrl_370;
  wire       [0:0]    _zz_ctrl_371;
  wire       [31:0]   _zz_ctrl_372;
  wire       [31:0]   _zz_ctrl_373;
  wire       [5:0]    _zz_ctrl_374;
  wire                _zz_ctrl_375;
  wire       [31:0]   _zz_ctrl_376;
  wire       [0:0]    _zz_ctrl_377;
  wire       [31:0]   _zz_ctrl_378;
  wire       [31:0]   _zz_ctrl_379;
  wire       [31:0]   _zz_ctrl_380;
  wire       [3:0]    _zz_ctrl_381;
  wire                _zz_ctrl_382;
  wire       [31:0]   _zz_ctrl_383;
  wire       [31:0]   _zz_ctrl_384;
  wire       [31:0]   _zz_ctrl_385;
  wire       [0:0]    _zz_ctrl_386;
  wire                _zz_ctrl_387;
  wire       [31:0]   _zz_ctrl_388;
  wire       [31:0]   _zz_ctrl_389;
  wire       [31:0]   _zz_ctrl_390;
  wire       [1:0]    _zz_ctrl_391;
  wire       [0:0]    _zz_ctrl_392;
  wire                _zz_ctrl_393;
  wire       [31:0]   _zz_ctrl_394;
  wire       [31:0]   _zz_ctrl_395;
  wire       [31:0]   _zz_ctrl_396;
  wire       [0:0]    _zz_ctrl_397;
  wire                _zz_ctrl_398;
  wire       [31:0]   _zz_ctrl_399;
  wire       [31:0]   _zz_ctrl_400;
  wire       [31:0]   _zz_ctrl_401;
  wire       [0:0]    _zz_ctrl_402;
  wire       [5:0]    _zz_ctrl_403;
  wire                _zz_ctrl_404;
  wire       [31:0]   _zz_ctrl_405;
  wire       [0:0]    _zz_ctrl_406;
  wire       [31:0]   _zz_ctrl_407;
  wire       [31:0]   _zz_ctrl_408;
  wire       [31:0]   _zz_ctrl_409;
  wire       [3:0]    _zz_ctrl_410;
  wire                _zz_ctrl_411;
  wire       [31:0]   _zz_ctrl_412;
  wire       [31:0]   _zz_ctrl_413;
  wire       [31:0]   _zz_ctrl_414;
  wire       [0:0]    _zz_ctrl_415;
  wire                _zz_ctrl_416;
  wire       [31:0]   _zz_ctrl_417;
  wire       [31:0]   _zz_ctrl_418;
  wire       [31:0]   _zz_ctrl_419;
  wire       [1:0]    _zz_ctrl_420;
  wire       [0:0]    _zz_ctrl_421;
  wire                _zz_ctrl_422;
  wire       [31:0]   _zz_ctrl_423;
  wire       [31:0]   _zz_ctrl_424;
  wire       [31:0]   _zz_ctrl_425;
  wire       [0:0]    _zz_ctrl_426;
  wire                _zz_ctrl_427;
  wire       [31:0]   _zz_ctrl_428;
  wire       [31:0]   _zz_ctrl_429;
  wire       [31:0]   _zz_ctrl_430;
  wire       [9:0]    _zz_ctrl_431;
  wire                _zz_ctrl_432;
  wire       [0:0]    _zz_ctrl_433;
  wire       [31:0]   _zz_ctrl_434;
  wire       [31:0]   _zz_ctrl_435;
  wire       [31:0]   _zz_ctrl_436;
  wire       [4:0]    _zz_ctrl_437;
  wire                _zz_ctrl_438;
  wire       [31:0]   _zz_ctrl_439;
  wire       [31:0]   _zz_ctrl_440;
  wire       [31:0]   _zz_ctrl_441;
  wire       [0:0]    _zz_ctrl_442;
  wire                _zz_ctrl_443;
  wire       [31:0]   _zz_ctrl_444;
  wire       [31:0]   _zz_ctrl_445;
  wire       [31:0]   _zz_ctrl_446;
  wire       [2:0]    _zz_ctrl_447;
  wire       [0:0]    _zz_ctrl_448;
  wire                _zz_ctrl_449;
  wire       [31:0]   _zz_ctrl_450;
  wire       [31:0]   _zz_ctrl_451;
  wire       [31:0]   _zz_ctrl_452;
  wire       [1:0]    _zz_ctrl_453;
  wire       [0:0]    _zz_ctrl_454;
  wire                _zz_ctrl_455;
  wire       [31:0]   _zz_ctrl_456;
  wire       [31:0]   _zz_ctrl_457;
  wire       [0:0]    _zz_ctrl_458;
  wire                _zz_ctrl_459;
  wire       [31:0]   _zz_ctrl_460;
  wire       [31:0]   _zz_ctrl_461;
  wire       [0:0]    _zz_ctrl_462;
  wire       [2:0]    _zz_ctrl_463;
  wire                _zz_ctrl_464;
  wire       [31:0]   _zz_ctrl_465;
  wire       [31:0]   _zz_ctrl_466;
  wire       [31:0]   _zz_ctrl_467;
  wire       [0:0]    _zz_ctrl_468;
  wire                _zz_ctrl_469;
  wire       [31:0]   _zz_ctrl_470;
  wire       [31:0]   _zz_ctrl_471;
  wire       [31:0]   _zz_ctrl_472;
  wire       [0:0]    _zz_ctrl_473;
  wire                _zz_ctrl_474;
  wire       [31:0]   _zz_ctrl_475;
  wire       [31:0]   _zz_ctrl_476;
  wire       [31:0]   _zz_ctrl_477;
  wire       [7:0]    _zz_ctrl_478;
  wire                _zz_ctrl_479;
  wire       [0:0]    _zz_ctrl_480;
  wire                _zz_ctrl_481;
  wire       [31:0]   _zz_ctrl_482;
  wire       [31:0]   _zz_ctrl_483;
  wire       [31:0]   _zz_ctrl_484;
  wire       [3:0]    _zz_ctrl_485;
  wire       [0:0]    _zz_ctrl_486;
  wire                _zz_ctrl_487;
  wire       [31:0]   _zz_ctrl_488;
  wire       [31:0]   _zz_ctrl_489;
  wire       [31:0]   _zz_ctrl_490;
  wire       [2:0]    _zz_ctrl_491;
  wire       [0:0]    _zz_ctrl_492;
  wire                _zz_ctrl_493;
  wire       [31:0]   _zz_ctrl_494;
  wire       [31:0]   _zz_ctrl_495;
  wire       [1:0]    _zz_ctrl_496;
  wire       [0:0]    _zz_ctrl_497;
  wire                _zz_ctrl_498;
  wire       [31:0]   _zz_ctrl_499;
  wire       [0:0]    _zz_ctrl_500;
  wire                _zz_ctrl_501;
  wire       [31:0]   _zz_ctrl_502;
  wire       [0:0]    _zz_ctrl_503;
  wire       [6:0]    _zz_ctrl_504;
  wire       [0:0]    _zz_ctrl_505;
  wire                _zz_ctrl_506;
  wire       [31:0]   _zz_ctrl_507;
  wire       [31:0]   _zz_ctrl_508;
  wire       [31:0]   _zz_ctrl_509;
  wire       [5:0]    _zz_ctrl_510;
  wire       [0:0]    _zz_ctrl_511;
  wire                _zz_ctrl_512;
  wire       [31:0]   _zz_ctrl_513;
  wire       [31:0]   _zz_ctrl_514;
  wire       [4:0]    _zz_ctrl_515;
  wire       [0:0]    _zz_ctrl_516;
  wire                _zz_ctrl_517;
  wire       [31:0]   _zz_ctrl_518;
  wire       [3:0]    _zz_ctrl_519;
  wire       [0:0]    _zz_ctrl_520;
  wire       [31:0]   _zz_ctrl_521;
  wire       [31:0]   _zz_ctrl_522;
  wire       [2:0]    _zz_ctrl_523;
  wire                _zz_ctrl_524;
  wire       [31:0]   _zz_ctrl_525;
  wire       [0:0]    _zz_ctrl_526;
  wire       [31:0]   _zz_ctrl_527;
  wire       [31:0]   _zz_ctrl_528;
  wire       [0:0]    _zz_ctrl_529;
  wire       [31:0]   _zz_ctrl_530;
  wire       [31:0]   _zz_ctrl_531;
  wire       [5:0]    _zz_ctrl_532;
  wire                _zz_ctrl_533;
  wire       [1:0]    _zz_ctrl_534;
  wire       [0:0]    _zz_ctrl_535;
  wire                _zz_ctrl_536;
  wire       [31:0]   _zz_ctrl_537;
  wire       [31:0]   _zz_ctrl_538;
  wire       [0:0]    _zz_ctrl_539;
  wire                _zz_ctrl_540;
  wire       [31:0]   _zz_ctrl_541;
  wire       [31:0]   _zz_ctrl_542;
  wire       [0:0]    _zz_ctrl_543;
  wire                _zz_ctrl_544;
  wire       [0:0]    _zz_ctrl_545;
  wire                _zz_ctrl_546;
  wire       [31:0]   _zz_ctrl_547;
  wire       [31:0]   _zz_ctrl_548;
  wire       [3:0]    _zz_ctrl_549;
  wire       [0:0]    _zz_ctrl_550;
  wire                _zz_ctrl_551;
  wire       [1:0]    _zz_ctrl_552;
  wire       [0:0]    _zz_ctrl_553;
  wire       [31:0]   _zz_ctrl_554;
  wire       [31:0]   _zz_ctrl_555;
  wire       [0:0]    _zz_ctrl_556;
  wire       [31:0]   _zz_ctrl_557;
  wire       [31:0]   _zz_ctrl_558;
  wire       [2:0]    _zz_ctrl_559;
  wire       [0:0]    _zz_ctrl_560;
  wire                _zz_ctrl_561;
  wire       [2:0]    _zz_ctrl_562;
  wire                _zz_ctrl_563;
  wire       [31:0]   _zz_ctrl_564;
  wire       [0:0]    _zz_ctrl_565;
  wire       [31:0]   _zz_ctrl_566;
  wire       [31:0]   _zz_ctrl_567;
  wire       [0:0]    _zz_ctrl_568;
  wire       [31:0]   _zz_ctrl_569;
  wire       [31:0]   _zz_ctrl_570;
  wire       [1:0]    _zz_ctrl_571;
  wire       [0:0]    _zz_ctrl_572;
  wire                _zz_ctrl_573;
  wire       [0:0]    _zz_ctrl_574;
  wire       [31:0]   _zz_ctrl_575;
  wire       [31:0]   _zz_ctrl_576;
  wire       [0:0]    _zz_ctrl_577;
  wire       [31:0]   _zz_ctrl_578;
  wire       [31:0]   _zz_ctrl_579;
  wire       [0:0]    _zz_ctrl_580;
  wire                _zz_ctrl_581;
  wire       [0:0]    _zz_ctrl_582;
  wire       [31:0]   _zz_ctrl_583;
  wire       [31:0]   _zz_ctrl_584;
  wire       [8:0]    _zz_ctrl_585;
  wire                _zz_ctrl_586;
  wire       [0:0]    _zz_ctrl_587;
  wire       [6:0]    _zz_ctrl_588;
  wire       [31:0]   _zz_ctrl_589;
  wire       [31:0]   _zz_ctrl_590;
  wire       [31:0]   _zz_ctrl_591;
  wire                _zz_ctrl_592;
  wire       [0:0]    _zz_ctrl_593;
  wire       [1:0]    _zz_ctrl_594;
  wire       [31:0]   _zz_fixInvalidInst;
  wire       [31:0]   _zz_fixInvalidInst_1;
  wire       [31:0]   _zz_fixInvalidInst_2;
  wire                _zz_fixInvalidInst_3;
  wire       [0:0]    _zz_fixInvalidInst_4;
  wire       [23:0]   _zz_fixInvalidInst_5;
  wire       [31:0]   _zz_fixInvalidInst_6;
  wire       [31:0]   _zz_fixInvalidInst_7;
  wire       [31:0]   _zz_fixInvalidInst_8;
  wire                _zz_fixInvalidInst_9;
  wire       [0:0]    _zz_fixInvalidInst_10;
  wire       [17:0]   _zz_fixInvalidInst_11;
  wire       [31:0]   _zz_fixInvalidInst_12;
  wire       [31:0]   _zz_fixInvalidInst_13;
  wire       [31:0]   _zz_fixInvalidInst_14;
  wire                _zz_fixInvalidInst_15;
  wire       [0:0]    _zz_fixInvalidInst_16;
  wire       [11:0]   _zz_fixInvalidInst_17;
  wire       [31:0]   _zz_fixInvalidInst_18;
  wire       [31:0]   _zz_fixInvalidInst_19;
  wire       [31:0]   _zz_fixInvalidInst_20;
  wire                _zz_fixInvalidInst_21;
  wire       [0:0]    _zz_fixInvalidInst_22;
  wire       [5:0]    _zz_fixInvalidInst_23;
  wire       [31:0]   _zz_fixInvalidInst_24;
  wire       [31:0]   _zz_fixInvalidInst_25;
  wire       [31:0]   _zz_fixInvalidInst_26;
  wire                _zz_fixInvalidInst_27;
  wire                _zz_fixInvalidInst_28;
  wire       [62:0]   ctrl;
  wire       [94:0]   fixDebug;
  wire       [95:0]   fixInvalidInst;

  assign _zz_ctrl = (inst_i & 32'h46409400);
  assign _zz_ctrl_1 = 32'h06400000;
  assign _zz_ctrl_2 = ((inst_i & 32'h46418000) == 32'h06408000);
  assign _zz_ctrl_3 = ((inst_i & 32'h66190000) == 32'h00090000);
  assign _zz_ctrl_4 = (|((inst_i & _zz_ctrl_5) == 32'h06000000));
  assign _zz_ctrl_6 = (|(_zz_ctrl_7 == _zz_ctrl_8));
  assign _zz_ctrl_9 = {(|_zz_ctrl_10),{(|_zz_ctrl_11),{_zz_ctrl_12,{_zz_ctrl_14,_zz_ctrl_17}}}};
  assign _zz_ctrl_5 = 32'h46400000;
  assign _zz_ctrl_7 = (inst_i & 32'h46408c00);
  assign _zz_ctrl_8 = 32'h06400000;
  assign _zz_ctrl_10 = ((inst_i & 32'h56000000) == 32'h04000000);
  assign _zz_ctrl_11 = ((inst_i & 32'h54008000) == 32'h10000000);
  assign _zz_ctrl_12 = (|((inst_i & _zz_ctrl_13) == 32'h10008000));
  assign _zz_ctrl_14 = (|(_zz_ctrl_15 == _zz_ctrl_16));
  assign _zz_ctrl_17 = {(|_zz_ctrl_18),{(|_zz_ctrl_19),{_zz_ctrl_20,{_zz_ctrl_33,_zz_ctrl_44}}}};
  assign _zz_ctrl_13 = 32'h54008000;
  assign _zz_ctrl_15 = (inst_i & 32'h46409400);
  assign _zz_ctrl_16 = 32'h06400400;
  assign _zz_ctrl_18 = ((inst_i & 32'h660c0000) == 32'h000c0000);
  assign _zz_ctrl_19 = ((inst_i & 32'h46408c00) == 32'h06400400);
  assign _zz_ctrl_20 = (|{(_zz_ctrl_21 == _zz_ctrl_22),{_zz_ctrl_23,{_zz_ctrl_25,_zz_ctrl_28}}});
  assign _zz_ctrl_33 = (|{_zz_ctrl_34,{_zz_ctrl_36,_zz_ctrl_39}});
  assign _zz_ctrl_44 = {(|_zz_ctrl_45),{(|_zz_ctrl_47),{_zz_ctrl_50,{_zz_ctrl_53,_zz_ctrl_60}}}};
  assign _zz_ctrl_21 = (inst_i & 32'h70000000);
  assign _zz_ctrl_22 = 32'h40000000;
  assign _zz_ctrl_23 = ((inst_i & _zz_ctrl_24) == 32'h10000000);
  assign _zz_ctrl_25 = (_zz_ctrl_26 == _zz_ctrl_27);
  assign _zz_ctrl_28 = {_zz_ctrl_29,_zz_ctrl_31};
  assign _zz_ctrl_34 = ((inst_i & _zz_ctrl_35) == 32'h40000000);
  assign _zz_ctrl_36 = (_zz_ctrl_37 == _zz_ctrl_38);
  assign _zz_ctrl_39 = {_zz_ctrl_40,_zz_ctrl_42};
  assign _zz_ctrl_45 = ((inst_i & _zz_ctrl_46) == 32'h06401800);
  assign _zz_ctrl_47 = (_zz_ctrl_48 == _zz_ctrl_49);
  assign _zz_ctrl_50 = (|_zz_ctrl_51);
  assign _zz_ctrl_53 = (|_zz_ctrl_54);
  assign _zz_ctrl_60 = {_zz_ctrl_61,{_zz_ctrl_69,_zz_ctrl_75}};
  assign _zz_ctrl_24 = 32'h70000000;
  assign _zz_ctrl_26 = (inst_i & 32'h68000000);
  assign _zz_ctrl_27 = 32'h40000000;
  assign _zz_ctrl_29 = ((inst_i & _zz_ctrl_30) == 32'h01000000);
  assign _zz_ctrl_31 = ((inst_i & _zz_ctrl_32) == 32'h00040000);
  assign _zz_ctrl_35 = 32'h70000000;
  assign _zz_ctrl_37 = (inst_i & 32'h70000000);
  assign _zz_ctrl_38 = 32'h10000000;
  assign _zz_ctrl_40 = ((inst_i & _zz_ctrl_41) == 32'h40000000);
  assign _zz_ctrl_42 = ((inst_i & _zz_ctrl_43) == 32'h000c0000);
  assign _zz_ctrl_46 = 32'h46409800;
  assign _zz_ctrl_48 = (inst_i & 32'h68000000);
  assign _zz_ctrl_49 = 32'h20000000;
  assign _zz_ctrl_51 = ((inst_i & _zz_ctrl_52) == 32'h01000000);
  assign _zz_ctrl_54 = {_zz_ctrl_55,{_zz_ctrl_56,_zz_ctrl_58}};
  assign _zz_ctrl_61 = (|{_zz_ctrl_62,_zz_ctrl_64});
  assign _zz_ctrl_69 = (|_zz_ctrl_70);
  assign _zz_ctrl_75 = {_zz_ctrl_76,{_zz_ctrl_79,_zz_ctrl_81}};
  assign _zz_ctrl_30 = 32'h61000000;
  assign _zz_ctrl_32 = 32'h664e0000;
  assign _zz_ctrl_41 = 32'h68000000;
  assign _zz_ctrl_43 = 32'h660c0000;
  assign _zz_ctrl_52 = 32'h53000000;
  assign _zz_ctrl_55 = ((inst_i & 32'h64000000) == 32'h44000000);
  assign _zz_ctrl_56 = ((inst_i & _zz_ctrl_57) == 32'h40000000);
  assign _zz_ctrl_58 = ((inst_i & _zz_ctrl_59) == 32'h40000000);
  assign _zz_ctrl_62 = ((inst_i & _zz_ctrl_63) == 32'h44000000);
  assign _zz_ctrl_64 = {(_zz_ctrl_65 == _zz_ctrl_66),(_zz_ctrl_67 == _zz_ctrl_68)};
  assign _zz_ctrl_70 = {(_zz_ctrl_71 == _zz_ctrl_72),(_zz_ctrl_73 == _zz_ctrl_74)};
  assign _zz_ctrl_76 = (|(_zz_ctrl_77 == _zz_ctrl_78));
  assign _zz_ctrl_79 = (|_zz_ctrl_80);
  assign _zz_ctrl_81 = {(|_zz_ctrl_82),{_zz_ctrl_83,{_zz_ctrl_85,_zz_ctrl_88}}};
  assign _zz_ctrl_57 = 32'h54000000;
  assign _zz_ctrl_59 = 32'h68000000;
  assign _zz_ctrl_63 = 32'h54000000;
  assign _zz_ctrl_65 = (inst_i & 32'h64000000);
  assign _zz_ctrl_66 = 32'h40000000;
  assign _zz_ctrl_67 = (inst_i & 32'h68000000);
  assign _zz_ctrl_68 = 32'h40000000;
  assign _zz_ctrl_71 = (inst_i & 32'h44000000);
  assign _zz_ctrl_72 = 32'h44000000;
  assign _zz_ctrl_73 = (inst_i & 32'h68000000);
  assign _zz_ctrl_74 = 32'h40000000;
  assign _zz_ctrl_77 = (inst_i & 32'h58000000);
  assign _zz_ctrl_78 = 32'h40000000;
  assign _zz_ctrl_80 = ((inst_i & 32'h70000000) == 32'h40000000);
  assign _zz_ctrl_82 = ((inst_i & 32'h40000000) == 32'h40000000);
  assign _zz_ctrl_83 = (|((inst_i & _zz_ctrl_84) == 32'h00200000));
  assign _zz_ctrl_85 = (|(_zz_ctrl_86 == _zz_ctrl_87));
  assign _zz_ctrl_88 = {(|_zz_ctrl_89),{(|_zz_ctrl_90),{_zz_ctrl_103,{_zz_ctrl_118,_zz_ctrl_139}}}};
  assign _zz_ctrl_84 = 32'h66280000;
  assign _zz_ctrl_86 = (inst_i & 32'h66280000);
  assign _zz_ctrl_87 = 32'h00200000;
  assign _zz_ctrl_89 = ((inst_i & 32'h66590000) == 32'h00080000);
  assign _zz_ctrl_90 = {(_zz_ctrl_91 == _zz_ctrl_92),{_zz_ctrl_93,{_zz_ctrl_95,_zz_ctrl_98}}};
  assign _zz_ctrl_103 = (|{_zz_ctrl_104,{_zz_ctrl_106,_zz_ctrl_109}});
  assign _zz_ctrl_118 = (|{_zz_ctrl_119,_zz_ctrl_122});
  assign _zz_ctrl_139 = {(|_zz_ctrl_140),{_zz_ctrl_155,{_zz_ctrl_156,_zz_ctrl_160}}};
  assign _zz_ctrl_91 = (inst_i & 32'h60000000);
  assign _zz_ctrl_92 = 32'h60000000;
  assign _zz_ctrl_93 = ((inst_i & _zz_ctrl_94) == 32'h58000000);
  assign _zz_ctrl_95 = (_zz_ctrl_96 == _zz_ctrl_97);
  assign _zz_ctrl_98 = {_zz_ctrl_99,_zz_ctrl_101};
  assign _zz_ctrl_104 = ((inst_i & _zz_ctrl_105) == 32'h60000000);
  assign _zz_ctrl_106 = (_zz_ctrl_107 == _zz_ctrl_108);
  assign _zz_ctrl_109 = {_zz_ctrl_110,{_zz_ctrl_112,_zz_ctrl_115}};
  assign _zz_ctrl_119 = (_zz_ctrl_120 == _zz_ctrl_121);
  assign _zz_ctrl_122 = {_zz_ctrl_123,{_zz_ctrl_125,_zz_ctrl_128}};
  assign _zz_ctrl_140 = {_zz_ctrl_141,{_zz_ctrl_143,_zz_ctrl_146}};
  assign _zz_ctrl_155 = 1'b0;
  assign _zz_ctrl_156 = (|_zz_ctrl_157);
  assign _zz_ctrl_160 = {_zz_ctrl_161,{_zz_ctrl_164,_zz_ctrl_176}};
  assign _zz_ctrl_94 = 32'h58000000;
  assign _zz_ctrl_96 = (inst_i & 32'h56000000);
  assign _zz_ctrl_97 = 32'h04000000;
  assign _zz_ctrl_99 = ((inst_i & _zz_ctrl_100) == 32'h02000000);
  assign _zz_ctrl_101 = ((inst_i & _zz_ctrl_102) == 32'h00100000);
  assign _zz_ctrl_105 = 32'h60000000;
  assign _zz_ctrl_107 = (inst_i & 32'h58000000);
  assign _zz_ctrl_108 = 32'h58000000;
  assign _zz_ctrl_110 = ((inst_i & _zz_ctrl_111) == 32'h04000000);
  assign _zz_ctrl_112 = (_zz_ctrl_113 == _zz_ctrl_114);
  assign _zz_ctrl_115 = (_zz_ctrl_116 == _zz_ctrl_117);
  assign _zz_ctrl_120 = (inst_i & 32'h70000000);
  assign _zz_ctrl_121 = 32'h40000000;
  assign _zz_ctrl_123 = ((inst_i & _zz_ctrl_124) == 32'h08000000);
  assign _zz_ctrl_125 = (_zz_ctrl_126 == _zz_ctrl_127);
  assign _zz_ctrl_128 = {_zz_ctrl_129,{_zz_ctrl_131,_zz_ctrl_134}};
  assign _zz_ctrl_141 = ((inst_i & _zz_ctrl_142) == 32'h10000000);
  assign _zz_ctrl_143 = (_zz_ctrl_144 == _zz_ctrl_145);
  assign _zz_ctrl_146 = {_zz_ctrl_147,{_zz_ctrl_149,_zz_ctrl_152}};
  assign _zz_ctrl_157 = (_zz_ctrl_158 == _zz_ctrl_159);
  assign _zz_ctrl_161 = (|_zz_ctrl_162);
  assign _zz_ctrl_164 = (|_zz_ctrl_165);
  assign _zz_ctrl_176 = {_zz_ctrl_177,{_zz_ctrl_196,_zz_ctrl_214}};
  assign _zz_ctrl_100 = 32'h67000000;
  assign _zz_ctrl_102 = 32'h721c0000;
  assign _zz_ctrl_111 = 32'h56000000;
  assign _zz_ctrl_113 = (inst_i & 32'h67000000);
  assign _zz_ctrl_114 = 32'h02000000;
  assign _zz_ctrl_116 = (inst_i & 32'h721c0000);
  assign _zz_ctrl_117 = 32'h00100000;
  assign _zz_ctrl_124 = 32'h68000000;
  assign _zz_ctrl_126 = (inst_i & 32'h6c000000);
  assign _zz_ctrl_127 = 32'h44000000;
  assign _zz_ctrl_129 = ((inst_i & _zz_ctrl_130) == 32'h01800000);
  assign _zz_ctrl_131 = (_zz_ctrl_132 == _zz_ctrl_133);
  assign _zz_ctrl_134 = {_zz_ctrl_135,_zz_ctrl_137};
  assign _zz_ctrl_142 = 32'h70000000;
  assign _zz_ctrl_144 = (inst_i & 32'h66400000);
  assign _zz_ctrl_145 = 32'h02400000;
  assign _zz_ctrl_147 = ((inst_i & _zz_ctrl_148) == 32'h00040000);
  assign _zz_ctrl_149 = (_zz_ctrl_150 == _zz_ctrl_151);
  assign _zz_ctrl_152 = (_zz_ctrl_153 == _zz_ctrl_154);
  assign _zz_ctrl_158 = (inst_i & 32'h70000000);
  assign _zz_ctrl_159 = 32'h10000000;
  assign _zz_ctrl_162 = ((inst_i & _zz_ctrl_163) == 32'h02000000);
  assign _zz_ctrl_165 = {_zz_ctrl_166,{_zz_ctrl_168,_zz_ctrl_171}};
  assign _zz_ctrl_177 = (|{_zz_ctrl_178,_zz_ctrl_181});
  assign _zz_ctrl_196 = (|_zz_ctrl_197);
  assign _zz_ctrl_214 = {_zz_ctrl_215,{_zz_ctrl_222,_zz_ctrl_226}};
  assign _zz_ctrl_130 = 32'h31800000;
  assign _zz_ctrl_132 = (inst_i & 32'h66210000);
  assign _zz_ctrl_133 = 32'h00010000;
  assign _zz_ctrl_135 = ((inst_i & _zz_ctrl_136) == 32'h00400000);
  assign _zz_ctrl_137 = ((inst_i & _zz_ctrl_138) == 32'h00008000);
  assign _zz_ctrl_148 = 32'h66140000;
  assign _zz_ctrl_150 = (inst_i & 32'h66190000);
  assign _zz_ctrl_151 = 32'h00010000;
  assign _zz_ctrl_153 = (inst_i & 32'h66608000);
  assign _zz_ctrl_154 = 32'h00008000;
  assign _zz_ctrl_163 = 32'h67000000;
  assign _zz_ctrl_166 = ((inst_i & _zz_ctrl_167) == 32'h00400000);
  assign _zz_ctrl_168 = (_zz_ctrl_169 == _zz_ctrl_170);
  assign _zz_ctrl_171 = {_zz_ctrl_172,_zz_ctrl_174};
  assign _zz_ctrl_178 = (_zz_ctrl_179 == _zz_ctrl_180);
  assign _zz_ctrl_181 = {_zz_ctrl_182,{_zz_ctrl_184,_zz_ctrl_187}};
  assign _zz_ctrl_197 = {_zz_ctrl_198,{_zz_ctrl_200,_zz_ctrl_203}};
  assign _zz_ctrl_215 = (|{_zz_ctrl_216,_zz_ctrl_219});
  assign _zz_ctrl_222 = (|_zz_ctrl_223);
  assign _zz_ctrl_226 = {_zz_ctrl_227,{_zz_ctrl_230,_zz_ctrl_236}};
  assign _zz_ctrl_136 = 32'h66480000;
  assign _zz_ctrl_138 = 32'h66508000;
  assign _zz_ctrl_167 = 32'h65400000;
  assign _zz_ctrl_169 = (inst_i & 32'h66280000);
  assign _zz_ctrl_170 = 32'h00080000;
  assign _zz_ctrl_172 = ((inst_i & _zz_ctrl_173) == 32'h02000000);
  assign _zz_ctrl_174 = ((inst_i & _zz_ctrl_175) == 32'h00020000);
  assign _zz_ctrl_179 = (inst_i & 32'h70000000);
  assign _zz_ctrl_180 = 32'h40000000;
  assign _zz_ctrl_182 = ((inst_i & _zz_ctrl_183) == 32'h10000000);
  assign _zz_ctrl_184 = (_zz_ctrl_185 == _zz_ctrl_186);
  assign _zz_ctrl_187 = {_zz_ctrl_188,{_zz_ctrl_190,_zz_ctrl_193}};
  assign _zz_ctrl_198 = ((inst_i & _zz_ctrl_199) == 32'h10000000);
  assign _zz_ctrl_200 = (_zz_ctrl_201 == _zz_ctrl_202);
  assign _zz_ctrl_203 = {_zz_ctrl_204,{_zz_ctrl_206,_zz_ctrl_209}};
  assign _zz_ctrl_216 = (_zz_ctrl_217 == _zz_ctrl_218);
  assign _zz_ctrl_219 = (_zz_ctrl_220 == _zz_ctrl_221);
  assign _zz_ctrl_223 = (_zz_ctrl_224 == _zz_ctrl_225);
  assign _zz_ctrl_227 = (|_zz_ctrl_228);
  assign _zz_ctrl_230 = (|_zz_ctrl_231);
  assign _zz_ctrl_236 = {_zz_ctrl_237,{_zz_ctrl_256,_zz_ctrl_274}};
  assign _zz_ctrl_173 = 32'h67800000;
  assign _zz_ctrl_175 = 32'h66220000;
  assign _zz_ctrl_183 = 32'h70000000;
  assign _zz_ctrl_185 = (inst_i & 32'h6c000000);
  assign _zz_ctrl_186 = 32'h44000000;
  assign _zz_ctrl_188 = ((inst_i & _zz_ctrl_189) == 32'h02000000);
  assign _zz_ctrl_190 = (_zz_ctrl_191 == _zz_ctrl_192);
  assign _zz_ctrl_193 = (_zz_ctrl_194 == _zz_ctrl_195);
  assign _zz_ctrl_199 = 32'h54000000;
  assign _zz_ctrl_201 = (inst_i & 32'h54008000);
  assign _zz_ctrl_202 = 32'h04008000;
  assign _zz_ctrl_204 = ((inst_i & _zz_ctrl_205) == 32'h04000000);
  assign _zz_ctrl_206 = (_zz_ctrl_207 == _zz_ctrl_208);
  assign _zz_ctrl_209 = {_zz_ctrl_210,_zz_ctrl_212};
  assign _zz_ctrl_217 = (inst_i & 32'h54400000);
  assign _zz_ctrl_218 = 32'h04400000;
  assign _zz_ctrl_220 = (inst_i & 32'h56000000);
  assign _zz_ctrl_221 = 32'h04000000;
  assign _zz_ctrl_224 = (inst_i & 32'h46410000);
  assign _zz_ctrl_225 = 32'h06410000;
  assign _zz_ctrl_228 = ((inst_i & _zz_ctrl_229) == 32'h00000400);
  assign _zz_ctrl_231 = {_zz_ctrl_232,_zz_ctrl_234};
  assign _zz_ctrl_237 = (|{_zz_ctrl_238,_zz_ctrl_241});
  assign _zz_ctrl_256 = (|_zz_ctrl_257);
  assign _zz_ctrl_274 = {_zz_ctrl_275,{_zz_ctrl_290,_zz_ctrl_296}};
  assign _zz_ctrl_189 = 32'h67000000;
  assign _zz_ctrl_191 = (inst_i & 32'h660c0000);
  assign _zz_ctrl_192 = 32'h000c0000;
  assign _zz_ctrl_194 = (inst_i & 32'h661c0000);
  assign _zz_ctrl_195 = 32'h00100000;
  assign _zz_ctrl_205 = 32'h56000000;
  assign _zz_ctrl_207 = (inst_i & 32'h54400000);
  assign _zz_ctrl_208 = 32'h04000000;
  assign _zz_ctrl_210 = ((inst_i & _zz_ctrl_211) == 32'h04000000);
  assign _zz_ctrl_212 = ((inst_i & _zz_ctrl_213) == 32'h04000000);
  assign _zz_ctrl_229 = 32'h66700400;
  assign _zz_ctrl_232 = ((inst_i & _zz_ctrl_233) == 32'h06410000);
  assign _zz_ctrl_234 = ((inst_i & _zz_ctrl_235) == 32'h00000000);
  assign _zz_ctrl_238 = (_zz_ctrl_239 == _zz_ctrl_240);
  assign _zz_ctrl_241 = {_zz_ctrl_242,{_zz_ctrl_244,_zz_ctrl_247}};
  assign _zz_ctrl_257 = {_zz_ctrl_258,{_zz_ctrl_260,_zz_ctrl_263}};
  assign _zz_ctrl_275 = (|{_zz_ctrl_276,_zz_ctrl_279});
  assign _zz_ctrl_290 = (|_zz_ctrl_291);
  assign _zz_ctrl_296 = {_zz_ctrl_297,{_zz_ctrl_312,_zz_ctrl_353}};
  assign _zz_ctrl_211 = 32'h54000800;
  assign _zz_ctrl_213 = 32'h54001000;
  assign _zz_ctrl_233 = 32'h46410000;
  assign _zz_ctrl_235 = 32'h66700400;
  assign _zz_ctrl_239 = (inst_i & 32'h71000000);
  assign _zz_ctrl_240 = 32'h01000000;
  assign _zz_ctrl_242 = ((inst_i & _zz_ctrl_243) == 32'h06410000);
  assign _zz_ctrl_244 = (_zz_ctrl_245 == _zz_ctrl_246);
  assign _zz_ctrl_247 = {_zz_ctrl_248,{_zz_ctrl_250,_zz_ctrl_253}};
  assign _zz_ctrl_258 = ((inst_i & _zz_ctrl_259) == 32'h01000000);
  assign _zz_ctrl_260 = (_zz_ctrl_261 == _zz_ctrl_262);
  assign _zz_ctrl_263 = {_zz_ctrl_264,{_zz_ctrl_266,_zz_ctrl_269}};
  assign _zz_ctrl_276 = (_zz_ctrl_277 == _zz_ctrl_278);
  assign _zz_ctrl_279 = {_zz_ctrl_280,{_zz_ctrl_282,_zz_ctrl_285}};
  assign _zz_ctrl_291 = {_zz_ctrl_292,_zz_ctrl_294};
  assign _zz_ctrl_297 = (|{_zz_ctrl_298,_zz_ctrl_301});
  assign _zz_ctrl_312 = (|_zz_ctrl_313);
  assign _zz_ctrl_353 = {_zz_ctrl_354,{_zz_ctrl_357,_zz_ctrl_369}};
  assign _zz_ctrl_243 = 32'h46410000;
  assign _zz_ctrl_245 = (inst_i & 32'h66400000);
  assign _zz_ctrl_246 = 32'h00400000;
  assign _zz_ctrl_248 = ((inst_i & _zz_ctrl_249) == 32'h00200000);
  assign _zz_ctrl_250 = (_zz_ctrl_251 == _zz_ctrl_252);
  assign _zz_ctrl_253 = (_zz_ctrl_254 == _zz_ctrl_255);
  assign _zz_ctrl_259 = 32'h51000000;
  assign _zz_ctrl_261 = (inst_i & 32'h46410000);
  assign _zz_ctrl_262 = 32'h06410000;
  assign _zz_ctrl_264 = ((inst_i & _zz_ctrl_265) == 32'h00400000);
  assign _zz_ctrl_266 = (_zz_ctrl_267 == _zz_ctrl_268);
  assign _zz_ctrl_269 = {_zz_ctrl_270,_zz_ctrl_272};
  assign _zz_ctrl_277 = (inst_i & 32'h68000000);
  assign _zz_ctrl_278 = 32'h20000000;
  assign _zz_ctrl_280 = ((inst_i & _zz_ctrl_281) == 32'h04000000);
  assign _zz_ctrl_282 = (_zz_ctrl_283 == _zz_ctrl_284);
  assign _zz_ctrl_285 = {_zz_ctrl_286,_zz_ctrl_288};
  assign _zz_ctrl_292 = ((inst_i & _zz_ctrl_293) == 32'h48000000);
  assign _zz_ctrl_294 = ((inst_i & _zz_ctrl_295) == 32'h20000000);
  assign _zz_ctrl_298 = (_zz_ctrl_299 == _zz_ctrl_300);
  assign _zz_ctrl_301 = {_zz_ctrl_302,{_zz_ctrl_304,_zz_ctrl_307}};
  assign _zz_ctrl_313 = {_zz_ctrl_314,{_zz_ctrl_316,_zz_ctrl_319}};
  assign _zz_ctrl_354 = (|_zz_ctrl_355);
  assign _zz_ctrl_357 = (|_zz_ctrl_358);
  assign _zz_ctrl_369 = {_zz_ctrl_370,{_zz_ctrl_402,_zz_ctrl_431}};
  assign _zz_ctrl_249 = 32'h66280000;
  assign _zz_ctrl_251 = (inst_i & 32'h660c0000);
  assign _zz_ctrl_252 = 32'h00040000;
  assign _zz_ctrl_254 = (inst_i & 32'h662c0000);
  assign _zz_ctrl_255 = 32'h00080000;
  assign _zz_ctrl_265 = 32'h66400000;
  assign _zz_ctrl_267 = (inst_i & 32'h66280000);
  assign _zz_ctrl_268 = 32'h00200000;
  assign _zz_ctrl_270 = ((inst_i & _zz_ctrl_271) == 32'h00040000);
  assign _zz_ctrl_272 = ((inst_i & _zz_ctrl_273) == 32'h00080000);
  assign _zz_ctrl_281 = 32'h54000000;
  assign _zz_ctrl_283 = (inst_i & 32'h54000000);
  assign _zz_ctrl_284 = 32'h10000000;
  assign _zz_ctrl_286 = ((inst_i & _zz_ctrl_287) == 32'h00080000);
  assign _zz_ctrl_288 = ((inst_i & _zz_ctrl_289) == 32'h00000000);
  assign _zz_ctrl_293 = 32'h48000000;
  assign _zz_ctrl_295 = 32'h28000000;
  assign _zz_ctrl_299 = (inst_i & 32'h48000000);
  assign _zz_ctrl_300 = 32'h48000000;
  assign _zz_ctrl_302 = ((inst_i & _zz_ctrl_303) == 32'h40000000);
  assign _zz_ctrl_304 = (_zz_ctrl_305 == _zz_ctrl_306);
  assign _zz_ctrl_307 = {_zz_ctrl_308,_zz_ctrl_310};
  assign _zz_ctrl_314 = ((inst_i & _zz_ctrl_315) == 32'h48000000);
  assign _zz_ctrl_316 = (_zz_ctrl_317 == _zz_ctrl_318);
  assign _zz_ctrl_319 = {_zz_ctrl_320,{_zz_ctrl_322,_zz_ctrl_325}};
  assign _zz_ctrl_355 = ((inst_i & _zz_ctrl_356) == 32'h08800000);
  assign _zz_ctrl_358 = {_zz_ctrl_359,{_zz_ctrl_361,_zz_ctrl_364}};
  assign _zz_ctrl_370 = (|{_zz_ctrl_371,_zz_ctrl_374});
  assign _zz_ctrl_402 = (|_zz_ctrl_403);
  assign _zz_ctrl_431 = {_zz_ctrl_432,{_zz_ctrl_462,_zz_ctrl_478}};
  assign _zz_ctrl_271 = 32'h660c0000;
  assign _zz_ctrl_273 = 32'h662c0000;
  assign _zz_ctrl_287 = 32'h72580000;
  assign _zz_ctrl_289 = 32'h72700000;
  assign _zz_ctrl_303 = 32'h50000000;
  assign _zz_ctrl_305 = (inst_i & 32'h1a000000);
  assign _zz_ctrl_306 = 32'h08000000;
  assign _zz_ctrl_308 = ((inst_i & _zz_ctrl_309) == 32'h08000000);
  assign _zz_ctrl_310 = ((inst_i & _zz_ctrl_311) == 32'h06000000);
  assign _zz_ctrl_315 = 32'h48000000;
  assign _zz_ctrl_317 = (inst_i & 32'h50000000);
  assign _zz_ctrl_318 = 32'h40000000;
  assign _zz_ctrl_320 = ((inst_i & _zz_ctrl_321) == 32'h00100000);
  assign _zz_ctrl_322 = (_zz_ctrl_323 == _zz_ctrl_324);
  assign _zz_ctrl_325 = {_zz_ctrl_326,{_zz_ctrl_328,_zz_ctrl_332}};
  assign _zz_ctrl_356 = 32'h5b800000;
  assign _zz_ctrl_359 = ((inst_i & _zz_ctrl_360) == 32'h00400000);
  assign _zz_ctrl_361 = (_zz_ctrl_362 == _zz_ctrl_363);
  assign _zz_ctrl_364 = {_zz_ctrl_365,_zz_ctrl_367};
  assign _zz_ctrl_371 = (_zz_ctrl_372 == _zz_ctrl_373);
  assign _zz_ctrl_374 = {_zz_ctrl_375,{_zz_ctrl_377,_zz_ctrl_381}};
  assign _zz_ctrl_403 = {_zz_ctrl_404,{_zz_ctrl_406,_zz_ctrl_410}};
  assign _zz_ctrl_432 = (|{_zz_ctrl_433,_zz_ctrl_437});
  assign _zz_ctrl_462 = (|_zz_ctrl_463);
  assign _zz_ctrl_478 = {_zz_ctrl_479,{_zz_ctrl_503,_zz_ctrl_532}};
  assign _zz_ctrl_309 = 32'h18800000;
  assign _zz_ctrl_311 = 32'h46400000;
  assign _zz_ctrl_321 = 32'h30100000;
  assign _zz_ctrl_323 = (inst_i & 32'h30800000);
  assign _zz_ctrl_324 = 32'h20000000;
  assign _zz_ctrl_326 = ((inst_i & _zz_ctrl_327) == 32'h04000000);
  assign _zz_ctrl_328 = (_zz_ctrl_329 == _zz_ctrl_331);
  assign _zz_ctrl_332 = {_zz_ctrl_333,{_zz_ctrl_337,_zz_ctrl_342}};
  assign _zz_ctrl_360 = 32'h64400000;
  assign _zz_ctrl_362 = (inst_i & 32'h66000000);
  assign _zz_ctrl_363 = 32'h02000000;
  assign _zz_ctrl_365 = ((inst_i & _zz_ctrl_366) == 32'h00100000);
  assign _zz_ctrl_367 = ((inst_i & _zz_ctrl_368) == 32'h00100000);
  assign _zz_ctrl_372 = (inst_i & 32'h70000000);
  assign _zz_ctrl_373 = 32'h40000000;
  assign _zz_ctrl_375 = ((inst_i & _zz_ctrl_376) == 32'h10000000);
  assign _zz_ctrl_377 = (_zz_ctrl_378 == _zz_ctrl_380);
  assign _zz_ctrl_381 = {_zz_ctrl_382,{_zz_ctrl_386,_zz_ctrl_391}};
  assign _zz_ctrl_404 = ((inst_i & _zz_ctrl_405) == 32'h60000000);
  assign _zz_ctrl_406 = (_zz_ctrl_407 == _zz_ctrl_409);
  assign _zz_ctrl_410 = {_zz_ctrl_411,{_zz_ctrl_415,_zz_ctrl_420}};
  assign _zz_ctrl_433 = (_zz_ctrl_434 == _zz_ctrl_436);
  assign _zz_ctrl_437 = {_zz_ctrl_438,{_zz_ctrl_442,_zz_ctrl_447}};
  assign _zz_ctrl_463 = {_zz_ctrl_464,{_zz_ctrl_468,_zz_ctrl_473}};
  assign _zz_ctrl_479 = (|{_zz_ctrl_480,_zz_ctrl_485});
  assign _zz_ctrl_503 = (|_zz_ctrl_504);
  assign _zz_ctrl_532 = {_zz_ctrl_533,{_zz_ctrl_543,_zz_ctrl_549}};
  assign _zz_ctrl_327 = 32'h16000000;
  assign _zz_ctrl_329 = (inst_i & _zz_ctrl_330);
  assign _zz_ctrl_331 = 32'h20000000;
  assign _zz_ctrl_333 = (_zz_ctrl_334 == _zz_ctrl_336);
  assign _zz_ctrl_337 = _zz_ctrl_338;
  assign _zz_ctrl_342 = {_zz_ctrl_343,_zz_ctrl_348};
  assign _zz_ctrl_366 = 32'h64180000;
  assign _zz_ctrl_368 = 32'h64140000;
  assign _zz_ctrl_376 = 32'h70000000;
  assign _zz_ctrl_378 = (inst_i & _zz_ctrl_379);
  assign _zz_ctrl_380 = 32'h40000000;
  assign _zz_ctrl_382 = (_zz_ctrl_383 == _zz_ctrl_385);
  assign _zz_ctrl_386 = _zz_ctrl_387;
  assign _zz_ctrl_391 = {_zz_ctrl_392,_zz_ctrl_397};
  assign _zz_ctrl_405 = 32'h60000000;
  assign _zz_ctrl_407 = (inst_i & _zz_ctrl_408);
  assign _zz_ctrl_409 = 32'h01000000;
  assign _zz_ctrl_411 = (_zz_ctrl_412 == _zz_ctrl_414);
  assign _zz_ctrl_415 = _zz_ctrl_416;
  assign _zz_ctrl_420 = {_zz_ctrl_421,_zz_ctrl_426};
  assign _zz_ctrl_434 = (inst_i & _zz_ctrl_435);
  assign _zz_ctrl_436 = 32'h10000000;
  assign _zz_ctrl_438 = (_zz_ctrl_439 == _zz_ctrl_441);
  assign _zz_ctrl_442 = _zz_ctrl_443;
  assign _zz_ctrl_447 = {_zz_ctrl_448,_zz_ctrl_453};
  assign _zz_ctrl_464 = (_zz_ctrl_465 == _zz_ctrl_467);
  assign _zz_ctrl_468 = _zz_ctrl_469;
  assign _zz_ctrl_473 = _zz_ctrl_474;
  assign _zz_ctrl_480 = _zz_ctrl_481;
  assign _zz_ctrl_485 = {_zz_ctrl_486,_zz_ctrl_491};
  assign _zz_ctrl_504 = {_zz_ctrl_505,_zz_ctrl_510};
  assign _zz_ctrl_533 = (|_zz_ctrl_534);
  assign _zz_ctrl_543 = _zz_ctrl_544;
  assign _zz_ctrl_549 = {_zz_ctrl_550,_zz_ctrl_559};
  assign _zz_ctrl_330 = 32'h32000000;
  assign _zz_ctrl_334 = (inst_i & _zz_ctrl_335);
  assign _zz_ctrl_336 = 32'h02000000;
  assign _zz_ctrl_338 = (_zz_ctrl_339 == _zz_ctrl_341);
  assign _zz_ctrl_343 = _zz_ctrl_344;
  assign _zz_ctrl_348 = _zz_ctrl_349;
  assign _zz_ctrl_379 = 32'h68000000;
  assign _zz_ctrl_383 = (inst_i & _zz_ctrl_384);
  assign _zz_ctrl_385 = 32'h06000000;
  assign _zz_ctrl_387 = (_zz_ctrl_388 == _zz_ctrl_390);
  assign _zz_ctrl_392 = _zz_ctrl_393;
  assign _zz_ctrl_397 = _zz_ctrl_398;
  assign _zz_ctrl_408 = 32'h41000000;
  assign _zz_ctrl_412 = (inst_i & _zz_ctrl_413);
  assign _zz_ctrl_414 = 32'h18000000;
  assign _zz_ctrl_416 = (_zz_ctrl_417 == _zz_ctrl_419);
  assign _zz_ctrl_421 = _zz_ctrl_422;
  assign _zz_ctrl_426 = _zz_ctrl_427;
  assign _zz_ctrl_435 = 32'h70000000;
  assign _zz_ctrl_439 = (inst_i & _zz_ctrl_440);
  assign _zz_ctrl_441 = 32'h00400000;
  assign _zz_ctrl_443 = (_zz_ctrl_444 == _zz_ctrl_446);
  assign _zz_ctrl_448 = _zz_ctrl_449;
  assign _zz_ctrl_453 = {_zz_ctrl_454,_zz_ctrl_458};
  assign _zz_ctrl_465 = (inst_i & _zz_ctrl_466);
  assign _zz_ctrl_467 = 32'h06000000;
  assign _zz_ctrl_469 = (_zz_ctrl_470 == _zz_ctrl_472);
  assign _zz_ctrl_474 = (_zz_ctrl_475 == _zz_ctrl_477);
  assign _zz_ctrl_481 = (_zz_ctrl_482 == _zz_ctrl_484);
  assign _zz_ctrl_486 = _zz_ctrl_487;
  assign _zz_ctrl_491 = {_zz_ctrl_492,_zz_ctrl_496};
  assign _zz_ctrl_505 = _zz_ctrl_506;
  assign _zz_ctrl_510 = {_zz_ctrl_511,_zz_ctrl_515};
  assign _zz_ctrl_534 = {_zz_ctrl_535,_zz_ctrl_539};
  assign _zz_ctrl_544 = (|_zz_ctrl_545);
  assign _zz_ctrl_550 = _zz_ctrl_551;
  assign _zz_ctrl_559 = {_zz_ctrl_560,_zz_ctrl_571};
  assign _zz_ctrl_335 = 32'h42400000;
  assign _zz_ctrl_339 = (inst_i & _zz_ctrl_340);
  assign _zz_ctrl_341 = 32'h00010000;
  assign _zz_ctrl_344 = (_zz_ctrl_345 == _zz_ctrl_347);
  assign _zz_ctrl_349 = (_zz_ctrl_350 == _zz_ctrl_352);
  assign _zz_ctrl_384 = 32'h46400000;
  assign _zz_ctrl_388 = (inst_i & _zz_ctrl_389);
  assign _zz_ctrl_390 = 32'h20000000;
  assign _zz_ctrl_393 = (_zz_ctrl_394 == _zz_ctrl_396);
  assign _zz_ctrl_398 = (_zz_ctrl_399 == _zz_ctrl_401);
  assign _zz_ctrl_413 = 32'h38000000;
  assign _zz_ctrl_417 = (inst_i & _zz_ctrl_418);
  assign _zz_ctrl_419 = 32'h04000000;
  assign _zz_ctrl_422 = (_zz_ctrl_423 == _zz_ctrl_425);
  assign _zz_ctrl_427 = (_zz_ctrl_428 == _zz_ctrl_430);
  assign _zz_ctrl_440 = 32'h64400000;
  assign _zz_ctrl_444 = (inst_i & _zz_ctrl_445);
  assign _zz_ctrl_446 = 32'h00100000;
  assign _zz_ctrl_449 = (_zz_ctrl_450 == _zz_ctrl_452);
  assign _zz_ctrl_454 = _zz_ctrl_455;
  assign _zz_ctrl_458 = _zz_ctrl_459;
  assign _zz_ctrl_466 = 32'h46400000;
  assign _zz_ctrl_470 = (inst_i & _zz_ctrl_471);
  assign _zz_ctrl_472 = 32'h20000000;
  assign _zz_ctrl_475 = (inst_i & _zz_ctrl_476);
  assign _zz_ctrl_477 = 32'h20000000;
  assign _zz_ctrl_482 = (inst_i & _zz_ctrl_483);
  assign _zz_ctrl_484 = 32'h20000000;
  assign _zz_ctrl_487 = (_zz_ctrl_488 == _zz_ctrl_490);
  assign _zz_ctrl_492 = _zz_ctrl_493;
  assign _zz_ctrl_496 = {_zz_ctrl_497,_zz_ctrl_500};
  assign _zz_ctrl_506 = (_zz_ctrl_507 == _zz_ctrl_509);
  assign _zz_ctrl_511 = _zz_ctrl_512;
  assign _zz_ctrl_515 = {_zz_ctrl_516,_zz_ctrl_519};
  assign _zz_ctrl_535 = _zz_ctrl_536;
  assign _zz_ctrl_539 = _zz_ctrl_540;
  assign _zz_ctrl_545 = _zz_ctrl_546;
  assign _zz_ctrl_551 = (|_zz_ctrl_552);
  assign _zz_ctrl_560 = _zz_ctrl_561;
  assign _zz_ctrl_571 = {_zz_ctrl_572,_zz_ctrl_580};
  assign _zz_ctrl_340 = 32'h30210000;
  assign _zz_ctrl_345 = (inst_i & _zz_ctrl_346);
  assign _zz_ctrl_347 = 32'h00400000;
  assign _zz_ctrl_350 = (inst_i & _zz_ctrl_351);
  assign _zz_ctrl_352 = 32'h00200000;
  assign _zz_ctrl_389 = 32'h70800000;
  assign _zz_ctrl_394 = (inst_i & _zz_ctrl_395);
  assign _zz_ctrl_396 = 32'h20000000;
  assign _zz_ctrl_399 = (inst_i & _zz_ctrl_400);
  assign _zz_ctrl_401 = 32'h000c0000;
  assign _zz_ctrl_418 = 32'h46000000;
  assign _zz_ctrl_423 = (inst_i & _zz_ctrl_424);
  assign _zz_ctrl_425 = 32'h00400000;
  assign _zz_ctrl_428 = (inst_i & _zz_ctrl_429);
  assign _zz_ctrl_430 = 32'h02000000;
  assign _zz_ctrl_445 = 32'h64100000;
  assign _zz_ctrl_450 = (inst_i & _zz_ctrl_451);
  assign _zz_ctrl_452 = 32'h02000000;
  assign _zz_ctrl_455 = (_zz_ctrl_456 == _zz_ctrl_457);
  assign _zz_ctrl_459 = (_zz_ctrl_460 == _zz_ctrl_461);
  assign _zz_ctrl_471 = 32'h70800000;
  assign _zz_ctrl_476 = 32'h72000000;
  assign _zz_ctrl_483 = 32'h68000000;
  assign _zz_ctrl_488 = (inst_i & _zz_ctrl_489);
  assign _zz_ctrl_490 = 32'h04000000;
  assign _zz_ctrl_493 = (_zz_ctrl_494 == _zz_ctrl_495);
  assign _zz_ctrl_497 = _zz_ctrl_498;
  assign _zz_ctrl_500 = _zz_ctrl_501;
  assign _zz_ctrl_507 = (inst_i & _zz_ctrl_508);
  assign _zz_ctrl_509 = 32'h20000000;
  assign _zz_ctrl_512 = (_zz_ctrl_513 == _zz_ctrl_514);
  assign _zz_ctrl_516 = _zz_ctrl_517;
  assign _zz_ctrl_519 = {_zz_ctrl_520,_zz_ctrl_523};
  assign _zz_ctrl_536 = (_zz_ctrl_537 == _zz_ctrl_538);
  assign _zz_ctrl_540 = (_zz_ctrl_541 == _zz_ctrl_542);
  assign _zz_ctrl_546 = (_zz_ctrl_547 == _zz_ctrl_548);
  assign _zz_ctrl_552 = {_zz_ctrl_553,_zz_ctrl_556};
  assign _zz_ctrl_561 = (|_zz_ctrl_562);
  assign _zz_ctrl_572 = _zz_ctrl_573;
  assign _zz_ctrl_580 = _zz_ctrl_581;
  assign _zz_ctrl_346 = 32'h64400000;
  assign _zz_ctrl_351 = 32'h30280000;
  assign _zz_ctrl_395 = 32'h72000000;
  assign _zz_ctrl_400 = 32'h460c0000;
  assign _zz_ctrl_424 = 32'h64400000;
  assign _zz_ctrl_429 = 32'h66000000;
  assign _zz_ctrl_451 = 32'h66000000;
  assign _zz_ctrl_456 = (inst_i & 32'h62410000);
  assign _zz_ctrl_457 = 32'h02410000;
  assign _zz_ctrl_460 = (inst_i & 32'h64280000);
  assign _zz_ctrl_461 = 32'h00200000;
  assign _zz_ctrl_489 = 32'h56000000;
  assign _zz_ctrl_494 = (inst_i & 32'h73000000);
  assign _zz_ctrl_495 = 32'h20000000;
  assign _zz_ctrl_498 = ((inst_i & _zz_ctrl_499) == 32'h20000000);
  assign _zz_ctrl_501 = ((inst_i & _zz_ctrl_502) == 32'h00000000);
  assign _zz_ctrl_508 = 32'h68000000;
  assign _zz_ctrl_513 = (inst_i & 32'h71000000);
  assign _zz_ctrl_514 = 32'h01000000;
  assign _zz_ctrl_517 = ((inst_i & _zz_ctrl_518) == 32'h00040000);
  assign _zz_ctrl_520 = (_zz_ctrl_521 == _zz_ctrl_522);
  assign _zz_ctrl_523 = {_zz_ctrl_524,{_zz_ctrl_526,_zz_ctrl_529}};
  assign _zz_ctrl_537 = (inst_i & 32'h73000000);
  assign _zz_ctrl_538 = 32'h20000000;
  assign _zz_ctrl_541 = (inst_i & 32'h71800000);
  assign _zz_ctrl_542 = 32'h20000000;
  assign _zz_ctrl_547 = (inst_i & 32'h62800000);
  assign _zz_ctrl_548 = 32'h22000000;
  assign _zz_ctrl_553 = (_zz_ctrl_554 == _zz_ctrl_555);
  assign _zz_ctrl_556 = (_zz_ctrl_557 == _zz_ctrl_558);
  assign _zz_ctrl_562 = {_zz_ctrl_563,{_zz_ctrl_565,_zz_ctrl_568}};
  assign _zz_ctrl_573 = (|{_zz_ctrl_574,_zz_ctrl_577});
  assign _zz_ctrl_581 = (|{_zz_ctrl_582,_zz_ctrl_585});
  assign _zz_ctrl_499 = 32'h71800000;
  assign _zz_ctrl_502 = 32'h72700000;
  assign _zz_ctrl_518 = 32'h66040000;
  assign _zz_ctrl_521 = (inst_i & 32'h73000000);
  assign _zz_ctrl_522 = 32'h20000000;
  assign _zz_ctrl_524 = ((inst_i & _zz_ctrl_525) == 32'h00400000);
  assign _zz_ctrl_526 = (_zz_ctrl_527 == _zz_ctrl_528);
  assign _zz_ctrl_529 = (_zz_ctrl_530 == _zz_ctrl_531);
  assign _zz_ctrl_554 = (inst_i & 32'h46400000);
  assign _zz_ctrl_555 = 32'h06000000;
  assign _zz_ctrl_557 = (inst_i & 32'h58800000);
  assign _zz_ctrl_558 = 32'h08000000;
  assign _zz_ctrl_563 = ((inst_i & _zz_ctrl_564) == 32'h20000000);
  assign _zz_ctrl_565 = (_zz_ctrl_566 == _zz_ctrl_567);
  assign _zz_ctrl_568 = (_zz_ctrl_569 == _zz_ctrl_570);
  assign _zz_ctrl_574 = (_zz_ctrl_575 == _zz_ctrl_576);
  assign _zz_ctrl_577 = (_zz_ctrl_578 == _zz_ctrl_579);
  assign _zz_ctrl_582 = (_zz_ctrl_583 == _zz_ctrl_584);
  assign _zz_ctrl_585 = {_zz_ctrl_586,{_zz_ctrl_587,_zz_ctrl_588}};
  assign _zz_ctrl_525 = 32'h66400000;
  assign _zz_ctrl_527 = (inst_i & 32'h71800000);
  assign _zz_ctrl_528 = 32'h20000000;
  assign _zz_ctrl_530 = (inst_i & 32'h66280000);
  assign _zz_ctrl_531 = 32'h00080000;
  assign _zz_ctrl_564 = 32'h68000000;
  assign _zz_ctrl_566 = (inst_i & 32'h60400000);
  assign _zz_ctrl_567 = 32'h20000000;
  assign _zz_ctrl_569 = (inst_i & 32'h46400000);
  assign _zz_ctrl_570 = 32'h06000000;
  assign _zz_ctrl_575 = (inst_i & 32'h6c000000);
  assign _zz_ctrl_576 = 32'h44000000;
  assign _zz_ctrl_578 = (inst_i & 32'h66700000);
  assign _zz_ctrl_579 = 32'h00000000;
  assign _zz_ctrl_583 = (inst_i & 32'h68000000);
  assign _zz_ctrl_584 = 32'h20000000;
  assign _zz_ctrl_586 = ((inst_i & 32'h70000000) == 32'h40000000);
  assign _zz_ctrl_587 = ((inst_i & 32'h46000000) == 32'h04000000);
  assign _zz_ctrl_588 = {((inst_i & 32'h6c000000) == 32'h44000000),{((inst_i & _zz_ctrl_589) == 32'h00400000),{(_zz_ctrl_590 == _zz_ctrl_591),{_zz_ctrl_592,{_zz_ctrl_593,_zz_ctrl_594}}}}};
  assign _zz_ctrl_589 = 32'h64400000;
  assign _zz_ctrl_590 = (inst_i & 32'h64100000);
  assign _zz_ctrl_591 = 32'h00100000;
  assign _zz_ctrl_592 = ((inst_i & 32'h66000000) == 32'h02000000);
  assign _zz_ctrl_593 = ((inst_i & 32'h73000000) == 32'h20000000);
  assign _zz_ctrl_594 = {((inst_i & 32'h64280000) == 32'h00200000),((inst_i & 32'h71800000) == 32'h20000000)};
  assign _zz_fixInvalidInst = 32'hdc000000;
  assign _zz_fixInvalidInst_1 = (inst_i & 32'hf6000000);
  assign _zz_fixInvalidInst_2 = 32'h14000000;
  assign _zz_fixInvalidInst_3 = ((inst_i & 32'hfe000000) == 32'h20000000);
  assign _zz_fixInvalidInst_4 = ((inst_i & 32'hfd800000) == 32'h28000000);
  assign _zz_fixInvalidInst_5 = {((inst_i & 32'hfe400000) == 32'h28000000),{((inst_i & 32'hfe800000) == 32'h28000000),{((inst_i & _zz_fixInvalidInst_6) == 32'h04000000),{(_zz_fixInvalidInst_7 == _zz_fixInvalidInst_8),{_zz_fixInvalidInst_9,{_zz_fixInvalidInst_10,_zz_fixInvalidInst_11}}}}}};
  assign _zz_fixInvalidInst_6 = 32'hff000000;
  assign _zz_fixInvalidInst_7 = (inst_i & 32'hff400000);
  assign _zz_fixInvalidInst_8 = 32'h2a400000;
  assign _zz_fixInvalidInst_9 = ((inst_i & 32'hff400000) == 32'h03400000);
  assign _zz_fixInvalidInst_10 = ((inst_i & 32'hfec00000) == 32'h02800000);
  assign _zz_fixInvalidInst_11 = {((inst_i & 32'hfec00000) == 32'h02400000),{((inst_i & 32'hfbc00000) == 32'h02000000),{((inst_i & _zz_fixInvalidInst_12) == 32'h00150000),{(_zz_fixInvalidInst_13 == _zz_fixInvalidInst_14),{_zz_fixInvalidInst_15,{_zz_fixInvalidInst_16,_zz_fixInvalidInst_17}}}}}};
  assign _zz_fixInvalidInst_12 = 32'hfffd0000;
  assign _zz_fixInvalidInst_13 = (inst_i & 32'hfff68000);
  assign _zz_fixInvalidInst_14 = 32'h00140000;
  assign _zz_fixInvalidInst_15 = ((inst_i & 32'hfff70000) == 32'h00140000);
  assign _zz_fixInvalidInst_16 = ((inst_i & 32'hfffe0000) == 32'h00200000);
  assign _zz_fixInvalidInst_17 = {((inst_i & 32'hfff38000) == 32'h00100000),{((inst_i & 32'hfffa8000) == 32'h00100000),{((inst_i & _zz_fixInvalidInst_18) == 32'h38720000),{(_zz_fixInvalidInst_19 == _zz_fixInvalidInst_20),{_zz_fixInvalidInst_21,{_zz_fixInvalidInst_22,_zz_fixInvalidInst_23}}}}}};
  assign _zz_fixInvalidInst_18 = 32'hffff0000;
  assign _zz_fixInvalidInst_19 = (inst_i & 32'hfffe8000);
  assign _zz_fixInvalidInst_20 = 32'h06488000;
  assign _zz_fixInvalidInst_21 = ((inst_i & 32'hfffe8000) == 32'h002a0000);
  assign _zz_fixInvalidInst_22 = ((inst_i & 32'hfffb8000) == 32'h00408000);
  assign _zz_fixInvalidInst_23 = {((inst_i & 32'hfff78000) == 32'h00408000),{((inst_i & 32'hffff0000) == 32'h00120000),{((inst_i & _zz_fixInvalidInst_24) == 32'h06483000),{(_zz_fixInvalidInst_25 == _zz_fixInvalidInst_26),{_zz_fixInvalidInst_27,_zz_fixInvalidInst_28}}}}};
  assign _zz_fixInvalidInst_24 = 32'hfffff800;
  assign _zz_fixInvalidInst_25 = (inst_i & 32'hfffff400);
  assign _zz_fixInvalidInst_26 = 32'h06483000;
  assign _zz_fixInvalidInst_27 = ((inst_i & 32'hfffff800) == 32'h06482800);
  assign _zz_fixInvalidInst_28 = ((inst_i & 32'hfffff800) == 32'h00006000);
  assign ctrl = {1'b0,{1'b0,{1'b0,{1'b0,{(|(_zz_ctrl == _zz_ctrl_1)),{(|_zz_ctrl_2),{(|_zz_ctrl_3),{_zz_ctrl_4,{_zz_ctrl_6,_zz_ctrl_9}}}}}}}}};
  assign fixDebug = {inst_i,ctrl};
  assign fixInvalidInst = {fixDebug,(! (|{((inst_i & 32'hf0000000) == 32'h50000000),{((inst_i & 32'hf0000000) == 32'h60000000),{((inst_i & _zz_fixInvalidInst) == 32'h4c000000),{(_zz_fixInvalidInst_1 == _zz_fixInvalidInst_2),{_zz_fixInvalidInst_3,{_zz_fixInvalidInst_4,_zz_fixInvalidInst_5}}}}}}))};
  assign is_o = fixInvalidInst;

endmodule
